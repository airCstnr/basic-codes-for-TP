
-- Variable
-- Une variable ne peut exister que dans un contexte séquentiel (= dans un process)

X := 1+2; -- X prend immédiatement la valeur 3 (sans pilote)

-- Eviter d’employer des variables, on leur préfèrera les signaux
-- Les variables sont principalement utilisées pour contenir les index des boucles
