
architecture simple of comparateur is
-- zone de déclaration (ici commentaire uniquement)
begin
-- zone de définition
egal <= ’1’ when a = b else ’0’; -- exemple d'architecture
end simple ;
