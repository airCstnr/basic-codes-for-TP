
-- Entité primaire de conception

-- En pratique, utilisez un fichier texte nom_entity.vhd pour chacune de vos entités nom_entity

entity nom_entity is
    -- port I/O
end entity nom_entity;
