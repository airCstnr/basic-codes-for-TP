
entity comparateur is
    port(
        a : in bit_vector(7 downto 0);
        b : in bit_vector(7 downto 0);
        egal : out bit);
end comparateur;
