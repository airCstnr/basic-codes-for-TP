
-- Architecture : définit les fonctionnalités et les relations temporelles

architecture nom_archi of nom_entité is
-- détailler le contenu
end architecture;
